`timescale 1ns / 1ps

module minesweeper_tb;

	/* == INPUTS == */
		reg			Clk;
		reg			Reset;
		reg			btnL;
		wire		btnL_Pulse;

	/* == OUTPUTS == */

	/* == PARAMETERS == */
		parameter x_size = 16;
		parameter y_size = 16;
		parameter x_coord_bits = 4;
		parameter y_coord_bits = 4;

	/* == LOCAL SIGNALS == */
		reg [(x_coord_bits - 1):0] x_coord;
		reg [(y_coord_bits - 1):0] y_coord;
		reg flag, open;
		wire [4:0] cell_val_board;
		wire [1:0] cell_val_cover;
		wire [(x_coord_bits + y_coord_bits - 1):0] num_mines;
		wire [31:0] rand, seed;
		wire game_over_wire;

	/* == INITIALIZE == */
		assign game_over_wire = (cell_val_cover[0] != 0) && (cell_val_board[4] != 0);

		initial begin
			Reset = 1;
			btnL = 0;
			x_coord = 0;
			y_coord = 0;
			flag = 0;
			open = 0;

			#20;
			Reset = 0;

			#103;

			#(16 * 16 * 20 * 2 + 100);

			#100;
			x_coord = 5'b00001;
			open = 1'b1;
			#20;
			open = 1'b0;
			#20;
		end

		initial begin
			Clk = 0;
			forever begin
				#10
				Clk = ~ Clk;
			end
		end

	/* == DESIGN == */
		debouncer #(.N_dc(7)) debouncer_L(
			.CLK(Clk), .RESET(Reset), .PB(btnL), .DPB( ), 
			.SCEN(btnL_Pulse), .MCEN( ), .CCEN( )
		);

		board board_arr(
			.clk(Clk), .reset(Reset),
			.x_coord(x_coord), .y_coord(y_coord),
			.cell_val(cell_val_board), .num_mines(num_mines),
			.seed(seed), .rand(rand),
			.is_init(), .init_x(), .init_y()
		);

		board_cover board_cover_arr(
			.clk(Clk), .reset(Reset),
			.flag(flag), .open(open),
			.x_coord(x_coord), .y_coord(y_coord),
			.cell_val(cell_val_cover)
		);

endmodule